library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library pll;
use pll.all;

entity telecran is
    port (
        -- FPGA
        i_clk_50: in std_logic;

        -- HDMI
        io_hdmi_i2c_scl       : inout std_logic;
        io_hdmi_i2c_sda       : inout std_logic;
        o_hdmi_tx_clk        : out std_logic;
        o_hdmi_tx_d          : out std_logic_vector(23 downto 0);
        o_hdmi_tx_de         : out std_logic;
        o_hdmi_tx_hs         : out std_logic;
        i_hdmi_tx_int        : in std_logic;
        o_hdmi_tx_vs         : out std_logic;

        -- KEYs
        i_rst_n : in std_logic;
		  
		-- LEDs
		o_leds : out std_logic_vector(9 downto 0);
		o_de10_leds : out std_logic_vector(7 downto 0);

		-- Coder
		i_left_ch_a : in std_logic;
		i_left_ch_b : in std_logic;
		i_left_pb : in std_logic;
		i_right_ch_a : in std_logic;
		i_right_ch_b : in std_logic;
		i_right_pb : in std_logic
    );
end entity telecran;

architecture rtl of telecran is
	component I2C_HDMI_Config 
		port (
			iCLK : in std_logic;
			iRST_N : in std_logic;
			I2C_SCLK : out std_logic;
			I2C_SDAT : inout std_logic;
			HDMI_TX_INT  : in std_logic
		);
	 end component;
	 
	component pll 
		port (
			refclk : in std_logic;
			rst : in std_logic;
			outclk_0 : out std_logic;
			locked : out std_logic
		);
	end component;

    constant h_res : natural := 720;
    constant v_res : natural := 480;
	 
	 signal h_val : natural;
	 signal v_val : natural;

	signal s_clk_27 : std_logic;
	signal s_rst_n : std_logic;	-- holds reset as long as pll is not locked
	
	signal a_prev, e : std_logic := '0';
begin
	o_leds <= (others => '0');
	o_de10_leds <= (others => '0');
	
	-- Frequency for HDMI is 27MHz generated by this PLL
	pll0 : component pll 
		port map (
			refclk => i_clk_50,
			rst => not(i_rst_n),
			outclk_0 => s_clk_27,
			locked => s_rst_n
		);

	-- Configures the ADV7513 for 480p
	I2C_HDMI_Config0 : component I2C_HDMI_Config 
		port map (
			iCLK => i_clk_50,
			iRST_N => i_rst_n,
			I2C_SCLK => io_hdmi_i2c_scl,
			I2C_SDAT => io_hdmi_i2c_sda,
			HDMI_TX_INT => i_hdmi_tx_int
	 );
	 
	 encodeur0 : component encodeur
	 generic map( MAX_COUNT =>v_res
	 );
		port map(
		  i_clk => i_clk_50,
        A    =>i_left_ch_a,
		  B    =>i_left_ch_b,
		  S 	 =>v_val
    );
	 
	 encodeur1 : component encodeur
	 generic map( MAX_COUNT =>h_res
	 );
		port map(
		  i_clk => i_clk_50,
        A    =>i_right_ch_a,
		  B    =>i_right_ch_b,
		  S 	 =>h_val
    );

	 
	 
end architecture rtl;
